LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY CW4 IS
	PORT ( SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	--wyświetlacze
	HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX4 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX5 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX6 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX7 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END CW4;

ARCHITECTURE strukturalna OF CW4 IS
	CONSTANT SPACJA: STD_LOGIC_VECTOR(2 DOWNTO 0):="000"; -- KOD SPACJI – uwaga na rodzaj ”” przy kompilacji

	--DEKLARACJA KOMPONENTÓW
	COMPONENT mux3bit8to1 -- muliptekser
		PORT ( 
			S, U0, U1, U2, U3, U4, U5,U6,U7: IN STD_LOGIC_VECTOR(2 DOWNTO 0); --WEKTOR STERUJĄCY I 8 wektorów INFORMACYJNYCH
			M : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
		);
	END COMPONENT;
	 
	COMPONENT char7seg -- transkoder
		PORT( 
			C : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			Display : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
			);
	END COMPONENT;
	 
	SIGNAL M0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL M1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL M2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL M3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL M4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL M5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL M6 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL M7 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	BEGIN
	-- KONKRETYZACJA UŻYCIA KOMPONENTÓW
	-- SW(17 DOWNTO 15) sterujący sygnal multipleksera
		-- DO WYKONANIA : KONKRETYZACJE KOLEJNYCH MULTIPLEKSERÓW UKŁADU
		MUX0: mux3bit8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),	SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA, M0);
		MUX1: mux3bit8to1 PORT MAP (SW(17 DOWNTO 15), SW(11 DOWNTO 9), SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA, SW(14 DOWNTO 12), M1);
		MUX2: mux3bit8to1 PORT MAP (SW(17 DOWNTO 15), SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA, SW(14 DOWNTO 12), SW(11 DOWNTO 9), M2);
		MUX3: mux3bit8to1 PORT MAP (SW(17 DOWNTO 15), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA, SW(14 DOWNTO 12), SW(11 DOWNTO 9), SW(8 DOWNTO 6), M3);
		MUX4: mux3bit8to1 PORT MAP (SW(17 DOWNTO 15), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA, SW(14 DOWNTO 12), SW(11 DOWNTO 9), SW(8 DOWNTO 6), SW(5 DOWNTO 3), M4);
		MUX5: mux3bit8to1 PORT MAP (SW(17 DOWNTO 15), SPACJA,SPACJA,SPACJA, SW(14 DOWNTO 12), SW(11 DOWNTO 9), SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),M5);
		MUX6: mux3bit8to1 PORT MAP (SW(17 DOWNTO 15), SPACJA,SPACJA, SW(14 DOWNTO 12), SW(11 DOWNTO 9), SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,M6);
		MUX7: mux3bit8to1 PORT MAP (SW(17 DOWNTO 15), SPACJA, SW(14 DOWNTO 12), SW(11 DOWNTO 9), SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,M7);
		-- DO WYKONANIA : KONKRETYZACJE KOLEJNYCH TRANSKODERÓW
		H0: char7seg PORT MAP (M0, HEX0);
		H1: char7seg PORT MAP (M1, HEX1);
		H2: char7seg PORT MAP (M2, HEX2);
		H3: char7seg PORT MAP (M3, HEX3);
		H4: char7seg PORT MAP (M4, HEX4);
		H5: char7seg PORT MAP (M5, HEX5);
		H6: char7seg PORT MAP (M6, HEX6);
		H7: char7seg PORT MAP (M7, HEX7);
	END strukturalna;